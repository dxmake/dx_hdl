module system_top (
);

system_wrapper system_wrapper_i (
);

endmodule
